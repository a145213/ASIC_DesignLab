// $Id: $
// File name:   test.sv
// Created:     11/16/2014
// Author:      Allen Chien
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: .
