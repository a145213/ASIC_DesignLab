library verilog;
use verilog.vl_types.all;
entity tb_flex_counter_8bit is
end tb_flex_counter_8bit;
