library verilog;
use verilog.vl_types.all;
entity tb_flex_counter_8bit_sv_unit is
end tb_flex_counter_8bit_sv_unit;
