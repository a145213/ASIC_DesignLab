// $Id: $
// File name:   adder_nbit.sv
// Created:     9/7/2014
// Author:      Allen Chien
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Creating a Parameterized Ripple Carry Adder Design

module adder_nbit
#(
  parameter BIT_WIDTH = 16
)
(
  input wire [(BIT_WIDTH - 1):0] a,
  input wire [(BIT_WIDTH - 1):0] b,
  input wire carry_in,
  output wire [(BIT_WIDTH - 1):0] sum,
  output wire overflow
);

wire [BIT_WIDTH:0] carrys;
genvar i;

assign carrys[0] = carry_in;
generate
  for(i = 0; i <= BIT_WIDTH - 1; i = i+1)
  begin
    adder_1bit IX (.a(a[i]), .b(b[i]), .carry_in(carrys[i]), .sum(sum[i]), .carry_out(carrys[i+1]));
  
  always @ (a)
  begin
    assert ((a[i] == 1'b0) || (a[i] == 1'b1))
      $info("input a correct");
    else 
      $error("input not correct");
  end

  always @ (b)
  begin
    assert ((b[i] == 1'b1) || (b[i] == 1'b0))
      $info("input b correct");
    else 
      $error("Input not correct");
  end

  always @ (a[i], b[i], carrys[i])
  begin
    assert (((a[i] + b[i] + carrys[i]) % 2) == sum[i])
      $info("output sum correct");
    else 
      $error("Output 's' of first 1 bit adder is not correct");
  end
  
  always @ (a[i], b[i], carry_in)
  begin
    assert ((((a[i] & b[i])|(carry_in & (a[i] ^ b[i]))) == carrys[i]))
      $info("carry correct");
    else
      $error("carry not correct");
  end
end
endgenerate

assign overflow = carrys[BIT_WIDTH];



endmodule